* adder circuit for tutorial

.model n nmos level=54
.model p pmos level=54

.subckt inv  in out
	mn1 out in gnd gnd n w=5.00u l=0.35u
	mp1 out in vdd vdd p w=10.00u l=0.35u
.ends

.subckt inv20  in out
	mn1 out in gnd gnd n w=20.00u l=0.35u
	mp1 out in vdd vdd p w=40.00u l=0.35u
.ends

.subckt xfer  gn gp d s
	mp1 d gp s vdd p w=10.00u l=0.35u
	mn1 d gn s gnd n w=5.00u l=0.35u
.ends

.subckt invr  in out
	mn1 out in gnd gnd n w=1.00u l=0.35u
	mp1 out in vdd vdd p w=2.00u l=0.35u
.ends

.subckt xor2  in1 in2 out
	mn1 out n3 n2 gnd n w=5.00u l=0.35u
	mp1 out n3 n4 vdd p w=10.00u l=0.35u
	x2  in2 n3 inv
	x3  n4 n2 inv 
	x4  n2 n4 n3 out xfer 
	x1  in1 n4 inv 
.ends

.subckt nor2  in1 in2 out
	mp1 n1 in1 vdd vdd p w=10.00u l=0.35u 
	mp2 out in2 n1 vdd p w=10.00u l=0.35u
	mn2 out in2 gnd gnd n w=5.00u l=0.35u
	mn1 out in1 gnd gnd n w=5.00u l=0.35u
.ends

.subckt addr  ain bin cout sum  cin
	x1  b  a  p  xor2
	x2 cin p sum xor2
	x3 bin bn inv20
	x4  bn b inv20
	x5 ain an inv20
	x6 an  a inv20
	x7 n1 n2 inv
	x8 b a k nor2
	x9 p k n1 nor2
	mn2 cout k gnd gnd n w=5.00u l=0.35u
	mp1 cout n2 vdd vdd p w=10.00u l=0.35u
	mn1 cout p cin gnd n w=5.00u l=0.35u
.ends

.subckt addr4 a_3 a_2 a_1 a_0 
+b_3 b_2 b_1 b_0 cin
+s_3 s_2 s_1 s_0 cout
	x1 a_3 b_3 cout s_3 n1 addr
	x2 a_2 b_2 n1 s_2 n2 addr
	x3 a_1 b_1 n2 s_1 n3 addr
	x4 a_0 b_0 n3 s_0 cin addr
.ends

.global vdd gnd
.print v(*)
vsu vdd gnd 3.3

.end
